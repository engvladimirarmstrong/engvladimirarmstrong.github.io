package sig_pkg;
  import uvm_pkg::*;
  `include "sig_item.svh"
  `include "sig_sequencer.svh"
  `include "sig_sequence.svh"
  `include "sig_driver.svh"
  `include "sig_monitor.svh"
  `include "sig_agent.svh"
  `include "sig_scoreboard.svh"
  `include "sig_model_env.svh"
  `include "sig_model_test.svh"
endpackage : sig_pkg
